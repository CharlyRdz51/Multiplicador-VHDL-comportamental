* Spice description of sum6bc_cougar
* Spice driver version -1218291655
* Date ( dd/mm/yyyy hh:mm:ss ):  9/02/2018 at 22:52:11

* INTERF a[0] a[1] a[2] a[3] a[4] a[5] b[0] b[1] b[2] b[3] b[4] b[5] cin 
* INTERF cout sum[0] sum[1] sum[2] sum[3] sum[4] sum[5] vdd vss 


.subckt sum6bc_cougar 248 251 175 167 143 187 249 250 135 69 227 188 233 156 
+ 228 196 81 44 15 110 255 226 
* NET 15 = sum[4]
* NET 23 = inv_x2_4_sig
* NET 24 = nao2o22_x1_sig
* NET 29 = not_aux21
* NET 31 = not_aux47
* NET 34 = na3_x1_sig
* NET 37 = no3_x1_sig
* NET 38 = noa22_x1_sig
* NET 41 = a2_x2_2_sig
* NET 44 = sum[3]
* NET 50 = na2_x1_2_sig
* NET 53 = mbk_buf_not_aux8
* NET 56 = no4_x1_sig
* NET 58 = a2_x2_sig
* NET 60 = o2_x2_sig
* NET 61 = not_b[2]
* NET 66 = xr2_x1_7_sig
* NET 69 = b[3]
* NET 81 = sum[2]
* NET 84 = mbk_buf_aux14
* NET 86 = na3_x1_4_sig
* NET 88 = inv_x2_2_sig
* NET 91 = aux16
* NET 95 = aux14
* NET 96 = not_aux14
* NET 98 = xr2_x1_6_sig
* NET 100 = not_a[2]
* NET 110 = sum[5]
* NET 114 = not_b[3]
* NET 115 = not_aux16
* NET 118 = not_a[3]
* NET 123 = inv_x2_5_sig
* NET 124 = not_aux17
* NET 125 = aux1
* NET 126 = not_aux49
* NET 132 = na4_x1_sig
* NET 135 = b[2]
* NET 136 = no2_x1_sig
* NET 141 = not_a[4]
* NET 143 = a[4]
* NET 145 = xr2_x1_9_sig
* NET 146 = nao22_x1_sig
* NET 152 = xr2_x1_8_sig
* NET 153 = na4_x1_2_sig
* NET 156 = cout
* NET 157 = inv_x2_3_sig
* NET 159 = not_aux8
* NET 160 = inv_x2_sig
* NET 162 = na2_x1_sig
* NET 163 = na3_x1_2_sig
* NET 164 = not_aux5
* NET 165 = not_b[0]
* NET 167 = a[3]
* NET 168 = aux6
* NET 175 = a[2]
* NET 180 = aux48
* NET 183 = aux0
* NET 187 = a[5]
* NET 188 = b[5]
* NET 189 = aux20
* NET 190 = ao22_x2_sig
* NET 196 = sum[1]
* NET 201 = not_cin
* NET 204 = aux13
* NET 208 = oa22_x2_sig
* NET 210 = not_b[1]
* NET 213 = mbk_buf_aux6
* NET 216 = xr2_x1_4_sig
* NET 220 = xr2_x1_5_sig
* NET 226 = vss
* NET 227 = b[4]
* NET 228 = sum[0]
* NET 233 = cin
* NET 234 = xr2_x1_sig
* NET 238 = xr2_x1_2_sig
* NET 241 = aux10
* NET 242 = not_aux10
* NET 244 = na2_x1_3_sig
* NET 245 = na3_x1_3_sig
* NET 246 = not_a[1]
* NET 247 = not_a[0]
* NET 248 = a[0]
* NET 249 = b[0]
* NET 250 = b[1]
* NET 251 = a[1]
* NET 254 = xr2_x1_3_sig
* NET 255 = vdd
Mtr_00478 244 250 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00477 255 251 244 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00476 246 251 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00475 255 249 245 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00474 245 251 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00473 245 248 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00472 252 251 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00471 255 250 253 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00470 254 252 256 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00469 256 250 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00468 256 253 254 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00467 255 251 256 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00466 241 237 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00465 255 248 237 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00464 237 249 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00463 242 241 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00462 240 241 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00461 255 254 243 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00460 238 240 239 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00459 239 254 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00458 239 243 238 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00457 255 241 239 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00456 247 248 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00455 232 249 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00454 255 233 236 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00453 234 232 235 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00452 235 233 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00451 235 236 234 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00450 255 249 235 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00449 230 248 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00448 255 234 231 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00447 228 230 229 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00446 229 234 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00445 229 231 228 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00444 255 248 229 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00443 219 251 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00442 255 250 222 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00441 220 219 176 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00440 176 250 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00439 176 222 220 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00438 255 251 176 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00437 201 233 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00436 217 213 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00435 255 220 218 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00434 216 217 174 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00433 174 220 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00432 174 218 216 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00431 255 213 174 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00430 210 250 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00429 172 216 197 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00428 172 201 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00427 255 238 172 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00426 197 233 172 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00425 196 197 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00424 255 242 204 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00423 204 244 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00422 204 201 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00421 255 207 208 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00420 173 210 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00419 173 242 207 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00418 207 246 173 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00417 255 192 190 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00416 192 189 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00415 255 187 171 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00414 171 188 192 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00413 178 188 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00412 255 187 184 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00411 180 178 170 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00410 170 187 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00409 170 184 180 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00408 255 188 170 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00407 183 191 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00406 255 187 191 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00405 191 188 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00404 168 165 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00403 255 247 168 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00402 160 168 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00401 255 246 166 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00400 164 166 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00399 255 247 166 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00398 166 165 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00397 213 169 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00396 255 168 169 255 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00395 255 158 159 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00394 158 210 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00393 255 160 161 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00392 161 246 158 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00391 144 180 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00390 255 146 147 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00389 145 144 148 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00388 148 146 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00387 148 147 145 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00386 255 180 148 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00385 255 162 163 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00384 163 213 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00383 163 233 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00382 162 210 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00381 255 246 162 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00380 255 155 156 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00379 155 153 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00378 255 190 154 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00377 154 183 155 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00376 157 183 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00375 149 180 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00374 255 189 150 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00373 152 149 151 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00372 151 189 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00371 151 150 152 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00370 255 180 151 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00369 141 143 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00368 165 249 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00367 108 141 136 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00366 255 135 108 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00365 255 136 132 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00364 132 208 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00363 255 163 132 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00362 132 245 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00361 255 141 125 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00360 125 128 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00359 255 227 128 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00358 123 125 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00357 255 124 146 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00356 106 126 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00355 146 123 106 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00354 255 118 153 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00353 153 126 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00352 255 157 153 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00351 153 124 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00350 105 115 113 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00349 255 114 105 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00348 126 113 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00347 102 145 109 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00346 102 167 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00345 255 152 102 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00344 109 118 102 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00343 110 109 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00342 96 95 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00341 88 204 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00340 100 175 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00339 255 164 90 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00338 89 159 95 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00337 90 88 89 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00336 189 87 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00335 255 125 87 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00334 87 86 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00333 99 175 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00332 255 135 101 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00331 98 99 97 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00330 97 135 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00329 97 101 98 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00328 255 175 97 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00327 91 93 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00326 94 175 92 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00325 94 135 255 255 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00324 255 175 94 255 tp L=1U W=14.5U AS=29P AD=29P PS=33U PD=33U 
Mtr_00323 92 135 93 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00322 93 95 94 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00321 84 85 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00320 255 95 85 255 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00319 80 98 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00318 255 84 83 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00317 81 80 82 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00316 82 84 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00315 82 83 81 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00314 255 98 82 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00313 115 91 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00312 255 114 86 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00311 86 115 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00310 86 124 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00309 58 76 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00308 255 96 76 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00307 76 61 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00306 61 135 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00305 255 143 52 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00304 54 53 55 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00303 55 61 56 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00302 52 164 54 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00301 59 96 77 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00300 255 61 59 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00299 60 77 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00298 53 73 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00297 255 159 73 255 tp L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00296 124 227 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00295 255 143 124 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00294 50 204 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00293 255 56 50 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00292 67 69 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00291 255 167 68 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00290 66 67 46 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00289 46 167 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00288 46 68 66 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00287 255 69 46 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00286 62 66 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00285 255 91 63 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00284 44 62 43 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00283 43 91 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00282 43 63 44 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00281 255 66 43 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00280 41 40 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00279 255 100 40 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00278 40 143 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00277 255 37 39 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00276 38 60 39 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00275 39 41 38 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00274 255 143 36 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00273 35 58 37 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00272 36 100 35 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00271 23 31 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00270 114 69 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00269 26 143 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00268 255 227 27 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00267 29 26 28 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00266 28 227 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00265 28 27 29 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00264 255 143 28 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00263 255 50 34 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00262 34 132 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00261 34 38 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00260 118 167 255 255 tp L=1U W=15U AS=30P AD=30P PS=34U PD=34U 
Mtr_00259 21 17 20 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00258 255 14 18 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00257 16 118 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00256 20 24 16 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00255 18 29 21 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00254 19 23 18 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00253 20 114 19 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00252 15 20 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00251 17 114 255 255 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00250 255 118 14 255 tp L=1U W=7U AS=14P AD=14P PS=18U PD=18U 
Mtr_00249 255 30 32 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00248 32 33 31 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00247 32 34 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00246 31 227 32 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00245 255 34 33 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00244 30 227 255 255 tp L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00243 24 29 25 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00242 25 114 255 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00241 22 69 24 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00240 255 31 22 255 tp L=1U W=20U AS=40P AD=40P PS=44U PD=44U 
Mtr_00239 226 250 209 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00238 209 251 244 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00237 226 251 246 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00236 226 248 211 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00235 211 249 212 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00234 212 251 245 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00233 253 250 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00232 226 251 252 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00231 224 252 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00230 254 253 224 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00229 225 251 254 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00228 226 250 225 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00227 237 249 195 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00226 226 237 241 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00225 195 248 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00224 226 241 242 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00223 243 254 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00222 226 241 240 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00221 200 240 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00220 238 243 200 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00219 199 241 238 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00218 226 254 199 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00217 226 248 247 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00216 236 233 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00215 226 249 232 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00214 186 232 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00213 234 236 186 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00212 194 249 234 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00211 226 233 194 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00210 231 234 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00209 226 248 230 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00208 182 230 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00207 228 231 182 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00206 181 248 228 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00205 226 234 181 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00204 222 250 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00203 226 251 219 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00202 223 219 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00201 220 222 223 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00200 221 251 220 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00199 226 250 221 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00198 226 233 201 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00197 218 220 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00196 226 213 217 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00195 215 217 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00194 216 218 215 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00193 214 213 216 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00192 226 220 214 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00191 226 250 210 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00190 203 216 197 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00189 226 233 203 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00188 198 201 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00187 197 238 198 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00186 226 197 196 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00185 226 201 205 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00184 205 242 202 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00183 202 244 204 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00182 208 207 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00181 226 210 207 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00180 206 242 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00179 207 246 206 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00178 192 187 193 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00177 193 188 192 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00176 226 189 193 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00175 190 192 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00174 184 187 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00173 226 188 178 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00172 179 178 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00171 180 184 179 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00170 177 188 180 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00169 226 187 177 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00168 191 188 185 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00167 226 191 183 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00166 185 187 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00165 226 165 142 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00164 142 247 168 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00163 226 168 160 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00162 226 166 164 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00161 139 246 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00160 140 165 139 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00159 166 247 140 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00158 226 169 213 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00157 169 168 226 226 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00156 158 160 130 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00155 130 246 158 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00154 226 210 130 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00153 159 158 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00152 147 146 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00151 226 180 144 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00150 111 144 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00149 145 147 111 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00148 112 180 145 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00147 226 146 112 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00146 226 233 133 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00145 133 162 134 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00144 134 213 163 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00143 226 210 129 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00142 129 246 162 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00141 155 190 122 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00140 122 183 155 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00139 226 153 122 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00138 156 155 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00137 226 183 157 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00136 150 189 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00135 226 180 149 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00134 116 149 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00133 152 150 116 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00132 117 180 152 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00131 226 189 117 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00130 226 143 141 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00129 226 249 165 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00128 136 135 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00127 226 141 136 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00126 226 245 138 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00125 138 136 137 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00124 137 208 131 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00123 131 163 132 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00122 128 227 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00121 107 141 125 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00120 226 128 107 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00119 226 125 123 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00118 127 126 146 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00117 146 123 127 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00116 127 124 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00115 226 124 121 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00114 121 118 119 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00113 119 126 120 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00112 120 157 153 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00111 126 113 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00110 113 114 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00109 226 115 113 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00108 104 145 109 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00107 226 118 104 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00106 103 167 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00105 109 152 103 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00104 226 109 110 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00103 226 95 96 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00102 226 204 88 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00101 226 175 100 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00100 226 88 95 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00099 95 164 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00098 95 159 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00097 87 86 72 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00096 226 87 189 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00095 72 125 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00094 101 135 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00093 226 175 99 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00092 78 99 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00091 98 101 78 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00090 79 175 98 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00089 226 135 79 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00088 226 93 91 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00087 226 135 74 226 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00086 74 175 226 226 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00085 93 135 75 226 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00084 75 175 226 226 tn L=1U W=9U AS=18P AD=18P PS=22U PD=22U 
Mtr_00083 74 95 93 226 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00082 226 85 84 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00081 85 95 226 226 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00080 83 84 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00079 226 98 80 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00078 64 80 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00077 81 83 64 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00076 65 98 81 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00075 226 84 65 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00074 226 91 115 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00073 226 124 71 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00072 71 114 70 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00071 70 115 86 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00070 76 61 57 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00069 226 76 58 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00068 57 96 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00067 226 135 61 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00066 56 143 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00065 226 61 56 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00064 226 164 56 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00063 56 53 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00062 60 77 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00061 77 61 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00060 226 96 77 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00059 226 73 53 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00058 73 159 226 226 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00057 226 227 49 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00056 49 143 124 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00055 226 204 51 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00054 51 56 50 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00053 68 167 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00052 226 69 67 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00051 48 67 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00050 66 68 48 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00049 47 69 66 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00048 226 167 47 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00047 63 91 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00046 226 66 62 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00045 42 62 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00044 44 63 42 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00043 45 66 44 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00042 226 91 45 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00041 40 143 13 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00040 226 40 41 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00039 13 100 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00038 226 60 12 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00037 12 41 38 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00036 38 37 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00035 226 100 37 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00034 37 143 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00033 37 58 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00032 226 31 23 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00031 226 69 114 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00030 27 227 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00029 226 143 26 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00028 6 26 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00027 29 27 6 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00026 7 143 29 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00025 226 227 7 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00024 226 38 11 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00023 11 50 10 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00022 10 132 34 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00021 226 167 118 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00020 226 114 17 226 tn L=1U W=4U AS=8P AD=8P PS=12U PD=12U 
Mtr_00019 14 118 226 226 tn L=1U W=3U AS=6P AD=6P PS=10U PD=10U 
Mtr_00018 4 29 2 226 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00017 2 114 20 226 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00016 20 17 3 226 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00015 3 23 4 226 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00014 226 118 4 226 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00013 1 14 226 226 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00012 20 24 1 226 tn L=1U W=6U AS=12P AD=12P PS=16U PD=16U 
Mtr_00011 226 20 15 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00010 226 34 9 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00009 9 30 31 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00008 31 33 8 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00007 8 227 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00006 226 227 30 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00005 33 34 226 226 tn L=1U W=5U AS=10P AD=10P PS=14U PD=14U 
Mtr_00004 226 31 5 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00003 5 69 226 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00002 24 29 5 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
Mtr_00001 5 114 24 226 tn L=1U W=10U AS=20P AD=20P PS=24U PD=24U 
C259 4 226 7.56e-15
C258 5 226 7.43e-15
C248 14 226 2.378e-14
C247 15 226 2.877e-14
C245 17 226 2.128e-14
C244 18 226 7.56e-15
C242 20 226 3.608e-14
C239 23 226 3.864e-14
C238 24 226 6.058e-14
C236 26 226 2.596e-14
C235 27 226 2.16e-14
C234 28 226 9.7e-15
C233 29 226 9.255e-14
C232 30 226 2.596e-14
C231 31 226 1.0773e-13
C230 32 226 7.76e-15
C229 33 226 2.16e-14
C228 34 226 5.561e-14
C225 37 226 5.407e-14
C224 38 226 5.697e-14
C223 39 226 6.05e-15
C222 40 226 1.8635e-14
C221 41 226 4.633e-14
C219 43 226 9.7e-15
C218 44 226 3.241e-14
C216 46 226 9.7e-15
C212 50 226 7.726e-14
C209 53 226 5.248e-14
C206 56 226 7.026e-14
C204 58 226 5.386e-14
C202 60 226 5.231e-14
C200 61 226 1.2246e-13
C199 62 226 2.596e-14
C198 63 226 2.16e-14
C195 66 226 7.195e-14
C194 67 226 2.596e-14
C193 68 226 2.16e-14
C192 69 226 1.6227e-13
C188 73 226 1.568e-14
C187 74 226 4.11e-15
C185 76 226 1.8635e-14
C184 77 226 1.8635e-14
C180 80 226 2.596e-14
C179 81 226 3.409e-14
C178 82 226 9.7e-15
C177 83 226 2.16e-14
C176 84 226 5.169e-14
C175 85 226 1.568e-14
C174 86 226 5.291e-14
C173 87 226 1.8635e-14
C172 88 226 5.064e-14
C169 91 226 1.2388e-13
C167 93 226 2.299e-14
C166 94 226 8.58e-15
C165 95 226 1.4248e-13
C164 96 226 9.534e-14
C163 97 226 9.7e-15
C162 98 226 1.3747e-13
C161 99 226 2.596e-14
C160 100 226 1.1929e-13
C159 101 226 2.16e-14
C158 102 226 7.43e-15
C150 109 226 2.445e-14
C149 110 226 6.523e-14
C146 113 226 1.8635e-14
C145 114 226 1.7562e-13
C144 115 226 7.885e-14
C141 118 226 1.7746e-13
C137 122 226 4.11e-15
C136 123 226 4.689e-14
C135 124 226 1.36e-13
C134 125 226 1.0926e-13
C133 126 226 8.547e-14
C132 127 226 4.11e-15
C131 128 226 1.662e-14
C129 130 226 4.11e-15
C127 132 226 8.168e-14
C124 135 226 1.8428e-13
C123 136 226 5.386e-14
C118 141 226 9.78e-14
C116 143 226 2.7541e-13
C114 144 226 2.596e-14
C113 145 226 5.245e-14
C112 146 226 8.473e-14
C111 147 226 2.16e-14
C110 148 226 9.7e-15
C109 149 226 2.596e-14
C108 150 226 2.16e-14
C107 151 226 9.7e-15
C106 152 226 6.085e-14
C105 153 226 5.749e-14
C103 155 226 1.853e-14
C102 156 226 5.063e-14
C101 157 226 5.784e-14
C100 158 226 1.853e-14
C99 159 226 1.0643e-13
C98 160 226 5.169e-14
C96 162 226 5.326e-14
C95 163 226 6.12e-14
C94 164 226 1.3819e-13
C93 165 226 8.558e-14
C92 166 226 2.605e-14
C91 167 226 2.324e-13
C90 168 226 1.2058e-13
C89 169 226 1.568e-14
C88 170 226 9.7e-15
C86 172 226 7.43e-15
C85 173 226 6.05e-15
C84 174 226 9.7e-15
C83 175 226 1.6725e-13
C81 176 226 9.7e-15
C79 178 226 2.596e-14
C77 180 226 1.0784e-13
C74 183 226 9.548e-14
C73 184 226 2.16e-14
C70 187 226 1.8246e-13
C69 188 226 9.868e-14
C68 189 226 1.1982e-13
C67 190 226 6.197e-14
C66 191 226 1.8635e-14
C65 192 226 1.853e-14
C64 193 226 4.11e-15
C61 196 226 8.155e-14
C60 197 226 2.445e-14
C56 201 226 9.2e-14
C53 204 226 1.2236e-13
C50 207 226 1.767e-14
C49 208 226 8.072e-14
C47 210 226 1.3187e-13
C44 213 226 1.1717e-13
C41 216 226 7.045e-14
C40 217 226 2.596e-14
C39 218 226 2.16e-14
C38 219 226 2.596e-14
C37 220 226 5.991e-14
C35 222 226 2.16e-14
C31 226 226 2.78936e-12
C30 227 226 2.7695e-13
C29 228 226 6.265e-14
C28 229 226 9.7e-15
C27 230 226 2.596e-14
C26 231 226 2.16e-14
C25 232 226 2.596e-14
C24 233 226 1.9823e-13
C23 234 226 5.751e-14
C22 235 226 9.7e-15
C21 236 226 2.16e-14
C20 237 226 1.8635e-14
C19 238 226 4.957e-14
C18 239 226 9.7e-15
C17 240 226 2.596e-14
C16 241 226 9.544e-14
C15 242 226 8.573e-14
C14 243 226 2.16e-14
C13 244 226 5.946e-14
C12 245 226 8.76e-14
C11 246 226 1.7549e-13
C10 247 226 8.865e-14
C9 248 226 1.9443e-13
C8 249 226 2.2162e-13
C7 250 226 2.1697e-13
C6 251 226 1.8534e-13
C5 252 226 2.596e-14
C4 253 226 2.16e-14
C3 254 226 8.991e-14
C2 255 226 2.89324e-12
C1 256 226 9.7e-15
.ends sum6bc_cougar

